// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_analog_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user analog project.
 *
 *-------------------------------------------------------------
 */

module user_analog_project_wrapper (
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    /* GPIOs.  There are 27 GPIOs, on either side of the analog.
     * These have the following mapping to the GPIO padframe pins
     * and memory-mapped registers, since the numbering remains the
     * same as caravel but skips over the analog I/O:
     *
     * io_in/out/oeb/in_3v3 [26:14]  <--->  mprj_io[37:25]
     * io_in/out/oeb/in_3v3 [13:0]   <--->  mprj_io[13:0]	
     *
     * When the GPIOs are configured by the Management SoC for
     * user use, they have three basic bidirectional controls:
     * in, out, and oeb (output enable, sense inverted).  For
     * analog projects, a 3.3V copy of the signal input is
     * available.  out and oeb must be 1.8V signals.
     */

    input  [`MPRJ_IO_PADS-`ANALOG_PADS-1:0] io_in,
    input  [`MPRJ_IO_PADS-`ANALOG_PADS-1:0] io_in_3v3,
    output [`MPRJ_IO_PADS-`ANALOG_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-`ANALOG_PADS-1:0] io_oeb,

    /* Analog (direct connection to GPIO pad---not for high voltage or
     * high frequency use).  The management SoC must turn off both
     * input and output buffers on these GPIOs to allow analog access.
     * These signals may drive a voltage up to the value of VDDIO
     * (3.3V typical, 5.5V maximum).
     * 
     * Note that analog I/O is not available on the 7 lowest-numbered
     * GPIO pads, and so the analog_io indexing is offset from the
     * GPIO indexing by 7, as follows:
     *
     * gpio_analog/noesd [17:7]  <--->  mprj_io[35:25]
     * gpio_analog/noesd [6:0]   <--->  mprj_io[13:7]	
     *
     */
    
    inout [`MPRJ_IO_PADS-`ANALOG_PADS-10:0] gpio_analog,
    inout [`MPRJ_IO_PADS-`ANALOG_PADS-10:0] gpio_noesd,

    /* Analog signals, direct through to pad.  These have no ESD at all,
     * so ESD protection is the responsibility of the designer.
     *
     * user_analog[10:0]  <--->  mprj_io[24:14]
     *
     */
    inout [`ANALOG_PADS-1:0] io_analog,

    /* Additional power supply ESD clamps, one per analog pad.  The
     * high side should be connected to a 3.3-5.5V power supply.
     * The low side should be connected to ground.
     *
     * clamp_high[2:0]   <--->  mprj_io[20:18]
     * clamp_low[2:0]    <--->  mprj_io[20:18]
     *
     */
    inout [2:0] io_clamp_high,
    inout [2:0] io_clamp_low,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_0();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_1();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_2();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_3();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_4();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_5();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_6();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_7();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_8();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_9();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_10();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_11();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_12();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_13();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_14();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_15();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_16();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_17();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_18();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_19();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_20();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_21();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_22();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_23();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_24();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_25();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_26();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_27();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_28();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_29();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_30();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_31();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_32();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_33();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_34();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_35();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_36();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_37();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_38();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_39();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_40();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_41();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_42();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_43();
M2M3_C_CDNS_641669455880 M2M3_C_CDNS_641669455880_44();

top_wrapper top_wrapper_0 (
//rram_LUT2 mprj (
//    `ifdef USE_POWER_PINS
//        .vdda1(vdda1),  // User area 1 3.3V power
//        .vdda2(vdda2),  // User area 2 3.3V power
//        .vssa1(vssa1),  // User area 1 analog ground
//        .vssa2(vssa2),  // User area 2 analog ground
//        .vccd1(vccd1),  // User area 1 1.8V power
//        .vccd2(vccd2),  // User area 2 1.8V power
//        .vssd1(vssd1),  // User area 1 digital ground
//        .vssd2(vssd2),  // User area 2 digital ground
//    `endif

    .vccd1(vccd1),  // User area 1 1.8V power
    .vdda1(vdda1),  // User area 1 1.8V power
    .vssd1(vssd1),  // User area 1 digital ground
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),

    // MGMT SoC Wishbone Slave

    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .wbs_sel_i(wbs_sel_i),
    .wbs_adr_i(wbs_adr_i),
    .wbs_dat_i(wbs_dat_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_dat_o(wbs_dat_o),

    // Logic Analyzer

    .la_data_in(la_data_in),
    .la_data_out(la_data_out),
    .la_oenb (la_oenb),

    // IO Pads
    .io_in (io_in),
    .io_in_3v3 (io_in_3v3),
    .io_out(io_out),
    .io_oeb(io_oeb),

    // GPIO-analog
    .gpio_analog(gpio_analog),
    .gpio_noesd(gpio_noesd),

    // Dedicated analog
    .io_analog(io_analog),
    .io_clamp_high(io_clamp_high),
    .io_clamp_low(io_clamp_low),

    // Clock
    .user_clock2(user_clock2),

    // IRQ
    .irq(user_irq)
);

endmodule	// user_analog_project_wrapper

`default_nettype wire
